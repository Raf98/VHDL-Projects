library verilog;
use verilog.vl_types.all;
entity ContadorAssinc3bits_vlg_vec_tst is
end ContadorAssinc3bits_vlg_vec_tst;
