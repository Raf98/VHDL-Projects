library verilog;
use verilog.vl_types.all;
entity Matrix_vlg_vec_tst is
end Matrix_vlg_vec_tst;
