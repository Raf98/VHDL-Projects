library verilog;
use verilog.vl_types.all;
entity FlipFlopJK_vlg_vec_tst is
end FlipFlopJK_vlg_vec_tst;
