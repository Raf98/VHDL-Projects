library verilog;
use verilog.vl_types.all;
entity Divisor_vlg_sample_tst is
    port(
        clock           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Divisor_vlg_sample_tst;
