library verilog;
use verilog.vl_types.all;
entity Contador4bits_vlg_vec_tst is
end Contador4bits_vlg_vec_tst;
