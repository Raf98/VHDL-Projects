library verilog;
use verilog.vl_types.all;
entity Functional_vlg_vec_tst is
end Functional_vlg_vec_tst;
