library verilog;
use verilog.vl_types.all;
entity bombaNova_vlg_vec_tst is
end bombaNova_vlg_vec_tst;
