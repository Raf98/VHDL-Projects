library verilog;
use verilog.vl_types.all;
entity Registrador1bit_vlg_vec_tst is
end Registrador1bit_vlg_vec_tst;
