library verilog;
use verilog.vl_types.all;
entity Contador3bits_vlg_vec_tst is
end Contador3bits_vlg_vec_tst;
